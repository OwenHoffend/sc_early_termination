module var_ET #(
    
)(

);

endmodule;